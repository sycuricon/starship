//VCS coverage exclude_file
`timescale 1ns / 10ps

`ifndef RESET_DELAY
  `define RESET_DELAY 15.7
`endif

`define SOC_TOP     Testbench.testHarness.ldut
`define TILE_TOP    `SOC_TOP.tile_prci_domain
`define MEM_TOP     Testbench.testHarness.mem.srams.mem
`define MEM_REG     `MEM_TOP.mem_ext

`ifdef TARGET_BOOM
  `define CPU_TOP   `TILE_TOP.tile_reset_domain_boom_tile
  `define PIPELINE  `CPU_TOP.core
  `define INTERRUPT `PIPELINE.io_interrupts_msip
`elsif TARGET_CVA6
  `define CPU_TOP   `TILE_TOP.tile_reset_domain_cva6_tile
  `define PIPELINE  `CPU_TOP.core.i_ariane.i_cva6
  `define INTERRUPT `PIPELINE.ipi_i
`elsif TARGET_XiangShan
  `define CPU_TOP   `TILE_TOP.tile_reset_domain_xiangshan_tile
  `define PIPELINE  `CPU_TOP.core.core.backend
  `define INTERRUPT `PIPELINE.io_externalInterrupt_msip
`else // TARGET_ROCKET
  `define CPU_TOP   `TILE_TOP.tile_reset_domain_tile
  `define PIPELINE  `CPU_TOP.core.core.backend
  `define INTERRUPT `PIPELINE.io_interrupts_msip
`endif

`ifdef COSIMULATION
  `define COVERAGE_PROBE Testbench.testHarness.ldut.io_covSum
  import "DPI-C" function int coverage_collector(
    input longint unsigned dut_cov
  );
  import "DPI-C" function void cosim_reinit(
      input string testcase,
      input reg verbose
  );
  import "DPI-C" function void cosim_set_tohost(input longint unsigned value);
`endif


module Testbench;
  
  reg clock = 1'b0;
  reg reset = 1'b1;

  wire interrupt;

  always #(`CLOCK_PERIOD/2.0) clock = ~clock;
  initial #(`RESET_DELAY) reset = 0;

  `ifdef VCS
    `ifdef COVERAGE_SUMMARY
      assign `SOC_TOP.metaReset = reset;
    `endif
  `endif

  initial begin
    `ifdef VCS
      `ifdef COVERAGE_SUMMARY
        force `INTERRUPT = interrupt;
      `endif
    `endif
  end 

  int unsigned rand_value;
  string testcase;
  string taintlog = "default";
  longint timer_result;
  
  reg [255:0] reason = "";
  reg failure = 1'b0;
  reg verbose = 1'b0;
  reg fuzzing = 1'b0;
  reg dump_wave = 1'b0;
  reg jtag_rbb_enable = 1'b0;
  reg [63:0] max_cycles = 0;
  reg [63:0] dump_start = 0;
  reg [63:0] trace_count = 0;
  reg [2047:0] fsdbfile = 0;
  reg [2047:0] vcdplusfile = 0;
  reg [2047:0] vcdfile = 0;

  int taint_fd;
  int event_fd;

  wire [63:0] tohost;
  wire printf_cond = verbose && !reset;
  wire uart_rx, uart_tx;

  initial begin
    void'($value$plusargs("max-cycles=%d", max_cycles));
    void'($value$plusargs("dump-start=%d", dump_start));
    void'($value$plusargs("jtag_rbb_enable=%d", jtag_rbb_enable));
    verbose = $test$plusargs("verbose");
    fuzzing = $test$plusargs("fuzzing");
    dump_wave = $test$plusargs("dump");

    // fixed for diffuzzRTL, CJ should not timeout
    max_cycles = 2000000000;

    // $urandom is seeded via cmdline (+ntb_random_seed in VCS) but that doesn't seed $random.
    rand_value = $urandom;
    rand_value = $random(rand_value);
    if (verbose) begin
      `ifdef VCS
        $fdisplay(32'h80000002, "testing $random %0x seed %d", rand_value, unsigned'($get_initial_random_seed));
      `endif
    end

    if (dump_wave) begin
      `ifdef DEBUG_FSDB
        `define WAVE_ON     $fsdbDumpon;
        `define WAVE_CLOSE  $fsdbDumpoff;
        $fsdbDumpfile({`TOP_DIR, "/wave/starship.fsdb"});
        $fsdbDumpvars(0, "+all");
      `elsif DEBUG_VCD
        `define WAVE_ON     $dumpon;
        `define WAVE_CLOSE  $dumpoff;
        $dumpfile({`TOP_DIR, "/wave/starship.vcd"});
        $dumpvars(0, Testbench);
      `else
        `define WAVE_ON     ;
        `define WAVE_CLOSE  ;
      `endif
    end

    if (dump_start == 0) begin
      // Start dumping before first clock edge to capture reset sequence in waveform
      if (dump_wave) begin
        `WAVE_ON
      end
    end
  end

  always @(negedge clock) begin
    if (!jtag_rbb_enable) begin
      trace_count = trace_count + 1;
      if (trace_count == dump_start) begin
        if (dump_wave) begin
          `WAVE_ON
        end
      end

      if (!reset) begin
        if (max_cycles > 0 && trace_count > max_cycles) begin
          reason = " (timeout)";
          failure = 1'b1;
        end

        if (failure) begin
          $fdisplay(32'h80000002, "*** FAILED ***%s after %d simulation cycles", reason, trace_count);
          trace_count = 0;
          failure = 0;
          `ifdef COSIMULATION
            if (fuzzing) begin
              $system("echo -e \"\033[31m[>] round timeout `date +%s.%3N` \033[0m\"");
              cosim_set_tohost(5);
              fuzz_manager();
            end
          `else
            if (dump_wave) begin
              `WAVE_CLOSE
            end
            $fatal;
          `endif
        end

        if (tohost & 1'b1) begin
          $fdisplay(32'h80000002, "*** PASSED *** Completed after %d simulation cycles", trace_count);
          trace_count = 0;
          `ifdef COSIMULATION
            if (fuzzing) begin
              $system("echo -e \"\033[31m[>] round finish `date +%s.%3N` \033[0m\"");
              fuzz_manager();
            end
          `else
            if (dump_wave) begin
              `WAVE_CLOSE
            end
            $system("echo -e \"\033[31m[>] vcs done `date +%s.%3N` \033[0m\"");
            `ifdef COVERAGE_SUMMARY
              $display("[CJ] coverage sum = %d", `COVERAGE_PROBE);
            `endif
            $finish;  
          `endif
        end
      end
    end
  end

  TestHarness testHarness(
    .clock(clock),
    .reset(reset),
    .io_uart_tx(),
    .io_uart_rx(1'b0)
  // .io_uart_tx(uart_tx),
  // .io_uart_rx(uart_rx)
  );

`ifdef COSIMULATION
  CJ rtlfuzz (
    .clock(clock),
    .reset(reset|jtag_rbb_enable),
    .tohost(tohost)
  );
`endif

  // tty #(115200, 0) u0_tty(
  //  .STX(uart_rx),
  //  .SRX(uart_tx),
  //  .reset(reset)
  // );

`ifdef COVERAGE_SUMMARY
  coverage_monitor mon(
    .clock(clock),
    .reset(reset),
    .cov(`COVERAGE_PROBE),
    .tohost(tohost),
    .interrupt(interrupt)
  );
`else
  assign interrupt = 0;
`endif

  task fuzz_manager;
  begin
    force clock = 0;
    #50;
    `ifdef COSIMULATION
      if (coverage_collector(`COVERAGE_PROBE)) begin
        reset = 1;
        $readmemh("./testcase.hex", `MEM_REG.ram);
        cosim_reinit("./testcase.elf", verbose);
        $system("echo -e \"\033[31m[>] round start `date +%s.%3N` \033[0m\"");
      end
    `endif
    release clock;
    #10 reset = 0;
  end
  endtask

endmodule


`define MAX_WAIT_CYCLE  1000

module coverage_monitor(
  input clock,
  input reset,
  input [29:0] cov,
  input [63:0] tohost,
  output interrupt
);

  reg [63:0] count = 0;
  reg [63:0] watch_dog = 0;
  reg [29:0] pre_cov = 0;

  always @(negedge clock) begin
    if (!reset) begin
      if (cov != pre_cov) begin
        pre_cov <= cov;
        count <= 0;
      end else begin
        count <= count + 1;
      end
      if (tohost & 1) begin
        count <= 0;
        watch_dog <= 0;
      end else begin
        watch_dog <= watch_dog + 1;
      end
    end else begin
      count <= 0;
      watch_dog <= 0;
    end
  end

  assign interrupt = (count >= (`MAX_WAIT_CYCLE * ((cov >> 19)+1) )) || (watch_dog >= 50000);
endmodule
